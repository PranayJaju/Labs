module AL3i(A, B, C, D, E, f);
    input A, B, C, D, E;
    output f;
    assign f=(~C&~D)|(A&~B&C&d);
endmodule 