module Q1a(A,lhs);
    input A;
    output lhs;
    assign lhs=~(~A);
endmodule