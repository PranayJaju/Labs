`timescale 1ns/1ns
`include "q1i.v"

module q1i_tb();
reg A, B, C;
wire Y;

q1i Q1i(A, B, C, Y);
initial
begin

    $dumpfile("q1i_tb.vcd");
    $dumpvars(0, q1i_tb);

    A=1'b0; B=1'b0; C=1'b0;
    #20;

    A=1'b0; B=1'b0; C=1'b1;
    #20;

    A=1'b0; B=1'b1; C=1'b0;
    #20;

    A=1'b0; B=1'b1; C=1'b1;
    #20;

    A=1'b1; B=1'b0; C=1'b0;
    #20;

    A=1'b1; B=1'b0; C=1'b1;
    #20;

    A=1'b1; B=1'b1; C=1'b0;
    #20;

    A=1'b1; B=1'b1; C=1'b1;
    #20;

    $display("Test complete");
end

endmodule